// Code your testbench here
// or browse Examples
module stim;
  wire [3:0]rdata;
  wire wfull, rempty;
  reg winc, rinc, rst, rclk, wclk;
  reg [3:0]wdata;
  
  CDC cdc1(wfull, rempty, rdata, winc, rinc, rst, rclk, wclk, wdata);
  initial $monitor(" At time=%0t, wdata=%h, wfull=%b, rempty=%b, rdata=%h, winc=%b, rst=%b",$time,wdata, wfull, rempty, rdata, winc, rst);
  
  //initial rempty=1, wfull=0;
  //initial rdata=4'b0000;
    initial begin
    $dumpfile("dump.vcd");
      $dumpvars(0);
  end
  initial begin 
    rclk=0; wclk=0; winc=1; rinc=1;
  end
  
  always 
    #5 wclk=~wclk;
  
  always
    #2 rclk=~rclk;
  
  always@(posedge wclk)
    begin
      winc <= (wfull==0)? 1:0;
    end

  
  initial begin
    rst=0; #30;
    wdata=4'b0110; #2;
    rst=1; #10;
    wdata=4'b0001; #10;
    wdata=4'b0010; #10;
    //$write("This is on ");
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
     wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    wdata=4'b0100; #10;
    wdata=4'b1000; #10;
    wdata=4'b0110; #10;
    wdata=4'b1100; #10;
    wdata=4'b0101; #10;
    wdata=4'b1010; #10;
    //$write("This is on fg ");
    wdata=4'b1111; #200;
    $finish;
  end
  
endmodule  