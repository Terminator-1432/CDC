`define WPTR_WIDTH 8
`define RPTR_WIDTH 8